//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "it"
//: property prefix = "_GG"
//: property title = "cubo.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] b;    //: /sn:0 {0}(#:160,177)(160,168)(160,168)(160,160){1}
//: {2}(162,158)(196,158){3}
//: {4}(200,158)(236,158){5}
//: {6}(198,156)(198,60)(591,60){7}
//: {8}(595,60)(698,60)(#:698,80){9}
//: {10}(593,62)(593,142)(635,142)(#:635,147){11}
//: {12}(158,158)(#:137,158){13}
reg [3:0] d;    //: /sn:0 {0}(#:697,290)(697,313)(606,313)(606,385){1}
//: {2}(608,387)(645,387)(#:645,366){3}
//: {4}(604,387)(221,387)(221,332){5}
//: {6}(223,330)(#:236,330){7}
//: {8}(219,330)(162,330){9}
//: {10}(158,330)(#:137,330){11}
//: {12}(160,332)(160,344)(160,344)(#:160,356){13}
reg [3:0] a;    //: /sn:0 {0}(#:236,105)(221,105){1}
//: {2}(219,103)(219,73)(602,73){3}
//: {4}(606,73)(648,73)(#:648,80){5}
//: {6}(604,75)(604,131)(701,131)(#:701,147){7}
//: {8}(217,105)(162,105){9}
//: {10}(160,103)(160,89)(160,89)(#:160,76){11}
//: {12}(158,105)(#:137,105){13}
reg [3:0] c;    //: /sn:0 {0}(#:137,275)(158,275){1}
//: {2}(162,275)(199,275){3}
//: {4}(203,275)(236,275){5}
//: {6}(201,277)(201,392)(597,392){7}
//: {8}(601,392)(689,392)(689,366){9}
//: {10}(599,390)(599,303)(638,303)(638,290){11}
//: {12}(160,273)(160,264)(160,264)(160,255){13}
wire [5:0] w6;    //: /sn:0 {0}(#:1183,162)(1183,207){1}
//: {2}(1185,209)(1250,209){3}
//: {4}(1181,209)(1145,209){5}
wire w7;    //: /sn:0 {0}(419,135)(450,135){1}
wire w16;    //: /sn:0 {0}(610,349)(590,349)(590,307){1}
//: {2}(590,303)(590,273)(610,273){3}
//: {4}(588,305)(575,305){5}
wire [3:0] w4;    //: /sn:0 {0}(#:763,91)(763,102){1}
//: {2}(761,104)(739,104){3}
//: {4}(#:763,106)(763,117)(807,117){5}
wire [4:0] w3;    //: /sn:0 {0}(#:941,133)(968,133){1}
//: {2}(972,133)(1026,133)(1026,194)(1036,194){3}
//: {4}(970,131)(970,100){5}
wire w0;    //: /sn:0 {0}(608,172)(588,172)(588,135){1}
//: {2}(588,131)(588,105)(610,105){3}
//: {4}(586,133)(575,133){5}
wire w1;    //: /sn:0 {0}(1404,185)(1423,185)(1423,143){1}
wire [5:0] w8;    //: /sn:0 {0}(#:1404,231)(1469,231)(1469,209){1}
wire [3:0] w17;    //: /sn:0 {0}(#:764,365)(764,350){1}
//: {2}(#:764,346)(764,327)(807,327){3}
//: {4}(762,348)(739,348){5}
wire [4:0] w10;    //: /sn:0 {0}(#:941,305)(968,305){1}
//: {2}(972,305)(1024,305)(1024,230)(1036,230){3}
//: {4}(970,303)(970,274){5}
wire [3:0] w13;    //: /sn:0 {0}(#:739,272)(761,272){1}
//: {2}(763,270)(#:763,263){3}
//: {4}(#:763,274)(763,289)(807,289){5}
wire w5;    //: /sn:0 {0}(450,307)(419,307){1}
wire [3:0] w9;    //: /sn:0 {0}(#:763,192)(763,173){1}
//: {2}(#:763,169)(763,155)(807,155){3}
//: {4}(761,171)(743,171){5}
//: enddecls

  //: LED g4 (a) @(160,69) /sn:0 /w:[ 11 ] /type:3
  //: joint g8 (d) @(160, 330) /w:[ 9 -1 10 12 ]
  //: joint g37 (w13) @(763, 272) /w:[ -1 2 1 4 ]
  sott4 g34 (.b(w9), .a(w4), .cout(w3));   //: @(808, 91) /sz:(132, 84) /sn:0 /p:[ Li0>3 Li1>5 Ro0<0 ]
  //: DIP g3 (d) @(99,330) /sn:0 /R:1 /w:[ 11 ] /st:0 /dn:1
  comparatore4 g13 (.a(c), .b(d), .c(w5));   //: @(237, 253) /sz:(181, 114) /sn:0 /p:[ Li0>5 Li1>7 Ro0<1 ]
  //: DIP g2 (c) @(99,275) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: DIP g1 (b) @(99,158) /sn:0 /R:1 /w:[ 13 ] /st:0 /dn:1
  mux4 g16 (.s(w16), .b(d), .a(c), .cout(w13));   //: @(611, 249) /sz:(127, 40) /sn:0 /p:[ Li0>3 Bi0>0 Bi1>11 Ro0<0 ]
  //: joint g11 (a) @(160, 105) /w:[ 9 10 12 -1 ]
  //: joint g10 (b) @(160, 158) /w:[ 2 -1 12 1 ]
  //: LED g28 (w4) @(763,84) /sn:0 /w:[ 0 ] /type:3
  inverter g19 (.a(w5), .cout(w16));   //: @(451, 284) /sz:(123, 48) /sn:0 /p:[ Li0>0 Ro0<5 ]
  //: joint g27 (b) @(593, 60) /w:[ 8 -1 7 10 ]
  //: joint g32 (c) @(599, 392) /w:[ 8 10 7 -1 ]
  //: joint g38 (w9) @(763, 171) /w:[ -1 2 4 1 ]
  //: LED g6 (c) @(160,248) /sn:0 /w:[ 13 ] /type:3
  //: joint g9 (c) @(160, 275) /w:[ 2 12 1 -1 ]
  //: LED g7 (d) @(160,363) /sn:0 /R:2 /w:[ 13 ] /type:3
  //: LED g31 (w17) @(764,372) /sn:0 /R:2 /w:[ 0 ] /type:3
  mux4 g15 (.b(a), .a(b), .s(w0), .cout(w9));   //: @(609, 148) /sz:(133, 40) /sn:0 /p:[ Ti0>7 Ti1>11 Li0>0 Ro0<5 ]
  //: joint g20 (w0) @(588, 133) /w:[ -1 2 4 1 ]
  //: joint g39 (w4) @(763, 104) /w:[ -1 1 2 4 ]
  //: joint g43 (w3) @(970, 133) /w:[ 2 4 1 -1 ]
  divisore g48 (.a(w6), .resto(w1), .cout(w8));   //: @(1251, 160) /sz:(152, 104) /sn:0 /p:[ Li0>3 Ro0<0 Ro1<0 ]
  //: LED g29 (w9) @(763,199) /sn:0 /R:2 /w:[ 0 ] /type:3
  mux4 g17 (.s(w16), .b(c), .a(d), .cout(w17));   //: @(611, 325) /sz:(127, 40) /sn:0 /p:[ Li0>0 Bi0>9 Bi1>3 Ro0<5 ]
  //: joint g25 (c) @(201, 275) /w:[ 4 -1 3 6 ]
  add5 g42 (.a(w3), .b(w10), .ris(w6));   //: @(1037, 166) /sz:(107, 85) /sn:0 /p:[ Li0>3 Li1>3 Ro0<5 ]
  mux4 g14 (.b(b), .a(a), .s(w0), .cout(w4));   //: @(611, 81) /sz:(127, 40) /sn:0 /p:[ Ti0>9 Ti1>5 Li0>3 Ro0<3 ]
  //: LED g5 (b) @(160,184) /sn:0 /R:2 /w:[ 0 ] /type:3
  //: joint g44 (w10) @(970, 305) /w:[ 2 4 1 -1 ]
  //: LED g47 (w1) @(1423,136) /sn:0 /w:[ 1 ] /type:0
  //: joint g36 (w17) @(764, 348) /w:[ -1 2 4 1 ]
  //: joint g21 (w16) @(590, 305) /w:[ -1 2 4 1 ]
  //: joint g24 (b) @(198, 158) /w:[ 4 6 3 -1 ]
  //: LED g41 (w3) @(970,93) /sn:0 /w:[ 5 ] /type:3
  //: joint g23 (a) @(219, 105) /w:[ 1 2 8 -1 ]
  //: LED g40 (w10) @(970,267) /sn:0 /w:[ 5 ] /type:3
  sott4 g35 (.b(w17), .a(w13), .cout(w10));   //: @(808, 263) /sz:(132, 84) /sn:0 /p:[ Li0>3 Li1>5 Ro0<0 ]
  //: DIP g0 (a) @(99,105) /sn:0 /R:1 /w:[ 13 ] /st:0 /dn:1
  //: joint g22 (d) @(221, 330) /w:[ 6 -1 8 5 ]
  //: joint g26 (a) @(604, 73) /w:[ 4 -1 3 6 ]
  //: LED g45 (w6) @(1183,155) /sn:0 /w:[ 0 ] /type:3
  //: joint g46 (w6) @(1183, 209) /w:[ 2 1 4 -1 ]
  comparatore4 g12 (.a(a), .b(b), .c(w7));   //: @(237, 81) /sz:(181, 114) /sn:0 /p:[ Li0>0 Li1>5 Ro0<0 ]
  inverter g18 (.a(w7), .cout(w0));   //: @(451, 112) /sz:(123, 48) /sn:0 /p:[ Li0>1 Ro0<5 ]
  //: joint g33 (d) @(606, 387) /w:[ 2 1 4 -1 ]
  //: LED g30 (w13) @(763,256) /sn:0 /w:[ 3 ] /type:3
  //: LED g49 (w8) @(1469,202) /sn:0 /w:[ 1 ] /type:3

endmodule
//: /netlistEnd

//: /netlistBegin add5
module add5(a, ris, b);
//: interface  /sz:(107, 85) /bd:[ Li0>a[4:0](28/85) Li1>b[4:0](64/85) Ro0<ris[5:0](43/85) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [4:0] b;    //: /sn:0 {0}(#:93,209)(196,209){1}
//: {2}(197,209)(357,209){3}
//: {4}(358,209)(443,209)(443,209)(505,209){5}
//: {6}(506,209)(562,209)(562,209)(658,209){7}
//: {8}(659,209)(861,209){9}
//: {10}(862,209)(876,209){11}
output [5:0] ris;    //: /sn:0 {0}(#:433,431)(433,484){1}
input [4:0] a;    //: /sn:0 {0}(#:93,143)(152,143){1}
//: {2}(153,143)(311,143){3}
//: {4}(312,143)(397,143)(397,143)(459,143){5}
//: {6}(460,143)(516,143)(516,143)(612,143){7}
//: {8}(613,143)(797,143){9}
//: {10}(798,143)(872,143){11}
wire w6;    //: /sn:0 {0}(160,321)(160,372)(410,372)(410,422){1}
wire w7;    //: /sn:0 {0}(896,302)(919,302)(919,400)(460,400)(460,422){1}
wire w14;    //: /sn:0 {0}(769,301)(723,301){1}
wire w16;    //: /sn:0 {0}(862,240)(862,213){1}
wire w4;    //: /sn:0 {0}(153,246)(153,157)(153,157)(153,147){1}
wire w15;    //: /sn:0 {0}(645,316)(645,358)(440,358)(440,422){1}
wire w0;    //: /sn:0 {0}(312,241)(312,155)(312,155)(312,147){1}
wire w3;    //: /sn:0 {0}(420,422)(420,358)(344,358)(344,318){1}
wire w21;    //: /sn:0 {0}(450,422)(450,382)(831,382)(831,320){1}
wire w1;    //: /sn:0 {0}(358,241)(358,188)(358,188)(358,213){1}
wire w8;    //: /sn:0 {0}(460,240)(460,147){1}
wire w18;    //: /sn:0 {0}(798,240)(798,147){1}
wire w17;    //: /sn:0 {0}(598,302)(570,302){1}
wire w12;    //: /sn:0 {0}(613,239)(613,147){1}
wire w2;    //: /sn:0 {0}(445,303)(435,303)(435,303)(422,303){1}
wire w11;    //: /sn:0 {0}(430,422)(430,340)(492,340)(492,317){1}
wire w10;    //: /sn:0 {0}(254,304)(297,304){1}
wire w13;    //: /sn:0 {0}(659,239)(659,213){1}
wire w5;    //: /sn:0 {0}(197,246)(197,190)(197,190)(197,213){1}
wire w9;    //: /sn:0 {0}(506,240)(506,213){1}
//: enddecls

  assign w1 = b[1]; //: TAP g8 @(358,207) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: IN g4 (a) @(91,143) /sn:0 /w:[ 0 ]
  full_adder g3 (.a(w12), .b(w13), .cin(w17), .s(w15), .cout(w14));   //: @(599, 240) /sz:(123, 75) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<0 Ro0<1 ]
  assign w13 = b[3]; //: TAP g13 @(659,207) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  full_adder g2 (.a(w8), .b(w9), .cin(w2), .s(w11), .cout(w17));   //: @(446, 241) /sz:(123, 75) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<1 ]
  full_adder g1 (.a(w0), .b(w1), .cin(w10), .s(w3), .cout(w2));   //: @(298, 242) /sz:(123, 75) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>1 Bo0<1 Ro0<1 ]
  assign w9 = b[2]; //: TAP g11 @(506,207) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  full_adder g16 (.a(w18), .b(w16), .cin(w14), .s(w21), .cout(w7));   //: @(770, 241) /sz:(125, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>0 Bo0<1 Ro0<0 ]
  assign w8 = a[2]; //: TAP g10 @(460,141) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign w4 = a[0]; //: TAP g6 @(153,141) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w0 = a[1]; //: TAP g9 @(312,141) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  assign w5 = b[0]; //: TAP g7 @(197,207) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: OUT g15 (ris) @(433,481) /sn:0 /R:3 /w:[ 1 ]
  assign w18 = a[4]; //: TAP g17 @(798,141) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1
  assign ris = {w7, w21, w15, w11, w3, w6}; //: CONCAT g14  @(435,427) /sn:0 /R:3 /w:[ 0 1 0 1 0 0 1 ] /dr:0 /tp:0 /drp:1
  //: IN g5 (b) @(91,209) /sn:0 /w:[ 0 ]
  half_adder g0 (.a(w4), .b(w5), .s(w6), .cout(w10));   //: @(130, 247) /sz:(123, 73) /sn:0 /p:[ Ti0>0 Ti1>0 Bo0<0 Ro0<0 ]
  assign w12 = a[3]; //: TAP g12 @(613,141) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w16 = b[4]; //: TAP g18 @(862,207) /sn:0 /R:1 /w:[ 1 9 10 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin divisore
module divisore(resto, cout, a);
//: interface  /sz:(152, 104) /bd:[ Li0>a[5:0](49/104) Ro0<resto(25/104) Ro1<cout[5:0](71/104) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output resto;    //: /sn:0 {0}(754,152)(754,195)(769,195){1}
//: {2}(773,195)(850,195){3}
//: {4}(771,197)(771,230){5}
supply1 w25;    //: /sn:0 {0}(694,258)(676,258)(676,222)(537,222){1}
//: {2}(533,222)(401,222){3}
//: {4}(397,222)(265,222){5}
//: {6}(261,222)(121,222){7}
//: {8}(117,222)(-26,222)(-26,256){9}
//: {10}(-24,258)(-4,258){11}
//: {12}(-28,258)(-53,258){13}
//: {14}(119,224)(119,258)(142,258){15}
//: {16}(263,224)(263,258)(278,258){17}
//: {18}(399,224)(399,258)(412,258){19}
//: {20}(535,224)(535,258)(554,258){21}
supply0 w2;    //: /sn:0 {0}(-46,158)(-46,215)(27,215)(27,230){1}
input [5:0] a;    //: /sn:0 {0}(#:94,148)(116,148){1}
//: {2}(117,148)(263,148){3}
//: {4}(264,148)(400,148){5}
//: {6}(401,148)(534,148){7}
//: {8}(535,148)(678,148){9}
//: {10}(679,148)(753,148){11}
//: {12}(754,148)(#:775,148){13}
output [5:0] cout;    //: /sn:0 {0}(#:397,507)(397,563){1}
wire w7;    //: /sn:0 {0}(402,501)(402,439)(464,439)(464,354){1}
wire w16;    //: /sn:0 {0}(173,230)(173,194)(119,194){1}
//: {2}(117,192)(117,152){3}
//: {4}(115,194)(73,194)(73,230){5}
wire w19;    //: /sn:0 {0}(48,354)(48,486)(372,486)(372,501){1}
wire w15;    //: /sn:0 {0}(382,501)(382,463)(194,463)(194,354){1}
wire w3;    //: /sn:0 {0}(412,501)(412,463)(606,463)(606,354){1}
wire w0;    //: /sn:0 {0}(631,230)(631,184)(677,184){1}
//: {2}(681,184)(725,184)(725,230){3}
//: {4}(679,182)(679,152){5}
wire w23;    //: /sn:0 {0}(746,354)(746,486)(422,486)(422,501){1}
wire w1;    //: /sn:0 {0}(585,230)(585,193)(537,193){1}
//: {2}(535,191)(535,152){3}
//: {4}(533,193)(489,193)(489,230){5}
wire w8;    //: /sn:0 {0}(443,230)(443,195)(403,195){1}
//: {2}(401,193)(401,152){3}
//: {4}(399,195)(355,195)(355,230){5}
wire w12;    //: /sn:0 {0}(309,230)(309,197)(266,197){1}
//: {2}(264,195)(264,152){3}
//: {4}(262,197)(219,197)(219,230){5}
wire w11;    //: /sn:0 {0}(392,501)(392,438)(330,438)(330,354){1}
//: enddecls

  //: VDD g8 (w25) @(-53,247) /sn:0 /R:1 /w:[ 13 ]
  shift1 g4 (.bit_succ(w16), .a(w12), .s(w25), .cout(w15));   //: @(143, 231) /sz:(100, 122) /sn:0 /p:[ Ti0>0 Ti1>5 Li0>15 Bo0<1 ]
  //: joint g13 (w25) @(535, 222) /w:[ 1 -1 2 20 ]
  shift1 g3 (.bit_succ(w12), .a(w8), .s(w25), .cout(w11));   //: @(279, 231) /sz:(100, 122) /sn:0 /p:[ Ti0>0 Ti1>5 Li0>17 Bo0<1 ]
  shift1 g2 (.bit_succ(w8), .a(w1), .s(w25), .cout(w7));   //: @(413, 231) /sz:(100, 122) /sn:0 /p:[ Ti0>0 Ti1>5 Li0>19 Bo0<1 ]
  shift1 g1 (.bit_succ(w1), .a(w0), .s(w25), .cout(w3));   //: @(555, 231) /sz:(100, 122) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>21 Bo0<1 ]
  //: joint g16 (resto) @(771, 195) /w:[ 2 -1 1 4 ]
  //: joint g11 (w25) @(263, 222) /w:[ 5 -1 6 16 ]
  //: joint g10 (w25) @(119, 222) /w:[ 7 -1 8 14 ]
  assign w12 = a[4]; //: TAP g28 @(264,146) /sn:0 /R:1 /w:[ 3 3 4 ] /ss:1
  //: joint g19 (w1) @(535, 193) /w:[ 1 2 4 -1 ]
  //: joint g27 (w12) @(264, 197) /w:[ 1 2 4 -1 ]
  shift1 g6 (.bit_succ(w0), .a(resto), .s(w25), .cout(w23));   //: @(695, 231) /sz:(100, 122) /sn:0 /p:[ Ti0>3 Ti1>5 Li0>0 Bo0<0 ]
  //: joint g9 (w25) @(-26, 258) /w:[ 10 9 12 -1 ]
  //: GROUND g7 (w2) @(-46,152) /sn:0 /R:2 /w:[ 0 ]
  assign w1 = a[2]; //: TAP g20 @(535,146) /sn:0 /R:1 /w:[ 3 7 8 ] /ss:1
  assign resto = a[0]; //: TAP g15 @(754,146) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  //: joint g17 (w0) @(679, 184) /w:[ 2 4 1 -1 ]
  //: joint g25 (w16) @(117, 194) /w:[ 1 2 4 -1 ]
  //: OUT g14 (resto) @(847,195) /sn:0 /w:[ 3 ]
  shift1 g5 (.bit_succ(w2), .a(w16), .s(w25), .cout(w19));   //: @(-3, 231) /sz:(100, 122) /sn:0 /p:[ Ti0>1 Ti1>5 Li0>11 Bo0<0 ]
  //: joint g21 (w8) @(401, 195) /w:[ 1 2 4 -1 ]
  assign cout = {w19, w15, w11, w7, w3, w23}; //: CONCAT g24  @(397,506) /sn:0 /R:3 /w:[ 0 1 0 0 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: OUT g23 (cout) @(397,560) /sn:0 /R:3 /w:[ 1 ]
  //: IN g0 (a) @(777,148) /sn:0 /R:2 /w:[ 13 ]
  assign w8 = a[3]; //: TAP g22 @(401,146) /sn:0 /R:1 /w:[ 3 5 6 ] /ss:1
  assign w16 = a[5]; //: TAP g26 @(117,146) /sn:0 /R:1 /w:[ 3 1 2 ] /ss:1
  assign w0 = a[1]; //: TAP g18 @(679,146) /sn:0 /R:1 /w:[ 5 9 10 ] /ss:1
  //: joint g12 (w25) @(399, 222) /w:[ 3 -1 4 18 ]

endmodule
//: /netlistEnd

//: /netlistBegin nand0
module nand0(a, b, cout);
//: interface  /sz:(93, 70) /bd:[ Li0>b(54/70) Li1>a(11/70) Ro0<cout(35/70) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(138,366)(226,366)(226,366)(168,366){1}
//: {2}(168,366)(239,366)(239,366)(249,366){3}
//: {4}(166,364)(166,213)(279,213){5}
supply0 w7;    //: /sn:0 {0}(263,498)(263,458){1}
supply1 w4;    //: /sn:0 {0}(259,112)(259,157){1}
//: {2}(261,159)(293,159)(293,205){3}
//: {4}(257,159)(230,159)(230,245){5}
input a;    //: /sn:0 {0}(138,253)(186,253){1}
//: {2}(190,253)(206,253)(206,253)(216,253){3}
//: {4}(188,255)(188,449)(249,449){5}
output cout;    //: /sn:0 {0}(263,358)(263,339){1}
//: {2}(265,337)(332,337){3}
//: {4}(263,335)(263,315){5}
//: {6}(265,313)(293,313)(293,222){7}
//: {8}(261,313)(230,313)(230,262){9}
wire w3;    //: /sn:0 {0}(263,441)(263,375){1}
//: enddecls

  //: IN g8 (a) @(136,253) /sn:0 /w:[ 0 ]
  //: joint g4 (cout) @(263, 313) /w:[ 6 -1 8 5 ]
  _GGNMOS #(2, 1) g3 (.Z(cout), .S(w3), .G(b));   //: @(257,366) /sn:0 /w:[ 0 1 3 ]
  //: joint g13 (cout) @(263, 337) /w:[ 2 4 -1 1 ]
  _GGNMOS #(2, 1) g2 (.Z(w3), .S(w7), .G(a));   //: @(257,449) /sn:0 /w:[ 0 1 5 ]
  _GGPMOS #(2, 1) g1 (.Z(cout), .S(w4), .G(b));   //: @(287,213) /sn:0 /w:[ 7 3 5 ]
  //: joint g11 (b) @(166, 366) /w:[ 2 4 1 -1 ]
  //: joint g10 (a) @(188, 253) /w:[ 2 -1 1 4 ]
  //: VDD g6 (w4) @(270,112) /sn:0 /w:[ 0 ]
  //: IN g9 (b) @(136,366) /sn:0 /w:[ 0 ]
  //: joint g7 (w4) @(259, 159) /w:[ 2 1 4 -1 ]
  //: GROUND g5 (w7) @(263,504) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) g0 (.Z(cout), .S(w4), .G(a));   //: @(224,253) /sn:0 /w:[ 9 5 3 ]
  //: OUT g12 (cout) @(329,337) /sn:0 /w:[ 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin and0
module and0(b, a, cout);
//: interface  /sz:(77, 48) /bd:[ Li0>a(8/48) Li1>b(36/48) Ro0<cout(23/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(29,221)(65,221){1}
input a;    //: /sn:0 {0}(30,178)(65,178){1}
output cout;    //: /sn:0 {0}(338,200)(316,200){1}
wire w2;    //: /sn:0 {0}(160,202)(191,202){1}
//: enddecls

  //: IN g4 (b) @(27,221) /sn:0 /w:[ 0 ]
  //: IN g3 (a) @(28,178) /sn:0 /w:[ 0 ]
  //: OUT g2 (cout) @(335,200) /sn:0 /w:[ 0 ]
  inverter g1 (.a(w2), .cout(cout));   //: @(192, 179) /sz:(123, 48) /sn:0 /p:[ Li0>1 Ro0<1 ]
  nand0 g0 (.b(b), .a(a), .cout(w2));   //: @(66, 167) /sz:(93, 70) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin and5
module and5(e, d, c, b, cout, a);
//: interface  /sz:(96, 94) /bd:[ Li0>e(81/94) Li1>d(64/94) Li2>c(44/94) Li3>b(27/94) Li4>a(8/94) Ro0<cout(44/94) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(255,222)(221,222)(221,222)(188,222){1}
input d;    //: /sn:0 {0}(255,257)(221,257)(221,257)(188,257){1}
input a;    //: /sn:0 {0}(188,203)(221,203)(221,203)(255,203){1}
output cout;    //: /sn:0 {0}(459,286)(497,286){1}
input c;    //: /sn:0 {0}(188,240)(220,240)(220,240)(255,240){1}
input e;    //: /sn:0 {0}(188,299)(285,299)(285,299)(380,299){1}
wire w4;    //: /sn:0 {0}(380,271)(354,271)(354,234)(339,234){1}
//: enddecls

  //: IN g4 (e) @(186,299) /sn:0 /w:[ 0 ]
  //: IN g3 (d) @(186,257) /sn:0 /w:[ 1 ]
  //: IN g2 (c) @(186,240) /sn:0 /w:[ 0 ]
  //: IN g1 (b) @(186,222) /sn:0 /w:[ 1 ]
  and0 g6 (.a(w4), .b(e), .cout(cout));   //: @(381, 263) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 ]
  //: OUT g7 (cout) @(494,286) /sn:0 /w:[ 1 ]
  and4 g5 (.d(d), .c(c), .b(b), .a(a), .cout(w4));   //: @(256, 186) /sz:(82, 82) /sn:0 /p:[ Li0>0 Li1>1 Li2>0 Li3>1 Ro0<1 ]
  //: IN g0 (a) @(186,203) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin full_add4
module full_add4(b, cout, a);
//: interface  /sz:(81, 103) /bd:[ Ti0>a[3:0](55/81) Ti1>b[3:0](29/81) Bo0<cout[4:0](44/81) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:199,195)(292,195){1}
//: {2}(293,195)(397,195){3}
//: {4}(398,195)(511,195){5}
//: {6}(512,195)(620,195){7}
//: {8}(621,195)(#:674,195){9}
supply1 w17;    //: /sn:0 {0}(701,296)(637,296){1}
input [3:0] a;    //: /sn:0 {0}(#:674,160)(589,160){1}
//: {2}(588,160)(484,160){3}
//: {4}(483,160)(370,160){5}
//: {6}(369,160)(262,160){7}
//: {8}(261,160)(203,160){9}
output [4:0] cout;    //: /sn:0 {0}(#:441,428)(441,479){1}
wire w6;    //: /sn:0 {0}(264,239)(264,172)(262,172)(262,164){1}
wire w7;    //: /sn:0 {0}(469,292)(414,292){1}
wire w14;    //: /sn:0 {0}(451,422)(451,375)(498,375)(498,319){1}
wire w19;    //: /sn:0 {0}(461,422)(461,398)(607,398)(607,321){1}
wire w4;    //: /sn:0 {0}(279,315)(279,383)(431,383)(431,422){1}
wire w15;    //: /sn:0 {0}(592,245)(592,172)(589,172)(589,164){1}
wire w3;    //: /sn:0 {0}(243,505)(243,525)(292,525)(292,401)(421,401)(421,422){1}
wire w0;    //: /sn:0 {0}(512,243)(512,199){1}
wire w1;    //: /sn:0 {0}(293,239)(293,199){1}
wire w8;    //: /sn:0 {0}(355,290)(309,290){1}
wire w12;    //: /sn:0 {0}(578,294)(528,294){1}
wire w2;    //: /sn:0 {0}(398,241)(398,199){1}
wire w11;    //: /sn:0 {0}(621,245)(621,199){1}
wire w10;    //: /sn:0 {0}(483,243)(483,172)(484,172)(484,164){1}
wire w13;    //: /sn:0 {0}(241,380)(241,288)(250,288){1}
wire w5;    //: /sn:0 {0}(369,241)(369,172)(370,172)(370,164){1}
wire w9;    //: /sn:0 {0}(441,422)(441,373)(384,373)(384,317){1}
//: enddecls

  assign w2 = b[2]; //: TAP g8 @(398,193) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  full_adder g4 (.b(w0), .a(w10), .cin(w12), .cout(w7), .s(w14));   //: @(470, 244) /sz:(57, 74) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  assign w15 = a[0]; //: TAP g13 @(589,158) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  full_adder g3 (.b(w2), .a(w5), .cin(w7), .cout(w8), .s(w9));   //: @(356, 242) /sz:(57, 74) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  full_adder g2 (.b(w1), .a(w6), .cin(w8), .cout(w13), .s(w4));   //: @(251, 240) /sz:(57, 74) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: IN g1 (b) @(676,195) /sn:0 /R:2 /w:[ 9 ]
  //: OUT g16 (cout) @(441,476) /sn:0 /R:3 /w:[ 1 ]
  assign w5 = a[2]; //: TAP g11 @(370,158) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  assign w6 = a[3]; //: TAP g10 @(262,158) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  assign w11 = b[0]; //: TAP g6 @(621,193) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  assign w1 = b[3]; //: TAP g9 @(293,193) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  assign w0 = b[1]; //: TAP g7 @(512,193) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  assign cout = {w3, w4, w9, w14, w19}; //: CONCAT g15  @(441,427) /sn:0 /R:3 /w:[ 0 1 1 0 0 0 ] /dr:1 /tp:0 /drp:1
  inverter g17 (.a(w13), .cout(w3));   //: @(216, 381) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  full_adder g5 (.b(w11), .a(w15), .cin(w17), .cout(w12), .s(w19));   //: @(579, 246) /sz:(57, 74) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: IN g0 (a) @(676,160) /sn:0 /R:2 /w:[ 0 ]
  assign w10 = a[1]; //: TAP g12 @(484,158) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  //: VDD g18 (w17) @(701,307) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin and3
module and3(c, b, cout, a);
//: interface  /sz:(75, 57) /bd:[ Li0>c(43/57) Li1>b(28/57) Li2>a(13/57) Ro0<cout(29/57) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(274,208)(339,208){1}
input a;    //: /sn:0 {0}(273,180)(339,180){1}
output cout;    //: /sn:0 {0}(604,210)(555,210){1}
input c;    //: /sn:0 {0}(271,242)(461,242)(461,223)(476,223){1}
wire w2;    //: /sn:0 {0}(476,195)(418,195){1}
//: enddecls

  and0 g4 (.a(w2), .b(c), .cout(cout));   //: @(477, 187) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>1 Ro0<1 ]
  //: IN g3 (c) @(269,242) /sn:0 /w:[ 0 ]
  //: IN g2 (b) @(272,208) /sn:0 /w:[ 0 ]
  and0 g1 (.a(a), .b(b), .cout(w2));   //: @(340, 172) /sz:(77, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 ]
  //: OUT g5 (cout) @(601,210) /sn:0 /w:[ 0 ]
  //: IN g0 (a) @(271,180) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin or0
module or0(b, a, cout);
//: interface  /sz:(57, 48) /bd:[ Li0>a(9/48) Li1>b(37/48) Ro0<cout(34/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(195,336)(221,336){1}
input a;    //: /sn:0 {0}(195,306)(221,306){1}
output cout;    //: /sn:0 {0}(451,329)(433,329){1}
wire w2;    //: /sn:0 {0}(285,331)(308,331){1}
//: enddecls

  //: IN g4 (b) @(193,336) /sn:0 /w:[ 0 ]
  //: IN g3 (a) @(193,306) /sn:0 /w:[ 0 ]
  //: OUT g2 (cout) @(448,329) /sn:0 /w:[ 0 ]
  nor0 g1 (.a(a), .b(b), .cout(w2));   //: @(222, 297) /sz:(62, 50) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  inverter g0 (.a(w2), .cout(cout));   //: @(309, 308) /sz:(123, 48) /sn:0 /p:[ Li0>1 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin sott4
module sott4(cout, b, a);
//: interface  /sz:(132, 84) /bd:[ Li0>a[3:0](26/84) Li1>b[3:0](64/84) Ro0<cout[4:0](42/84) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:114,245)(114,290){1}
input [3:0] a;    //: /sn:0 {0}(#:230,313)(230,401){1}
output [4:0] cout;    //: /sn:0 {0}(#:219,596)(219,506){1}
wire [3:0] w0;    //: /sn:0 {0}(#:119,343)(119,367)(204,367)(204,401){1}
//: enddecls

  //: OUT g4 (cout) @(219,593) /sn:0 /R:3 /w:[ 0 ]
  full_add4 g3 (.b(w0), .a(a), .cout(cout));   //: @(175, 402) /sz:(81, 103) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]
  complemento g2 (.b(b), .cout(w0));   //: @(19, 291) /sz:(194, 51) /sn:0 /p:[ Ti0>1 Bo0<0 ]
  //: IN g1 (b) @(114,243) /sn:0 /R:3 /w:[ 0 ]
  //: IN g0 (a) @(230,311) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin half_adder
module half_adder(a, cout, s, b);
//: interface  /sz:(64, 73) /bd:[ Ti0>a(45/64) Ti1>b(19/64) Lo0<cout(52/73) Bo0<s(38/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(95,57)(65,57)(65,154){1}
//: {2}(67,156)(165,156){3}
//: {4}(63,156)(52,156){5}
output s;    //: /sn:0 {0}(271,41)(204,41)(204,41)(196,41){1}
input a;    //: /sn:0 {0}(48,29)(99,29)(99,29)(81,29){1}
//: {2}(81,29)(103,29)(103,29)(95,29){3}
//: {4}(79,31)(79,128)(165,128){5}
output cout;    //: /sn:0 {0}(271,143)(244,143){1}
//: enddecls

  //: IN g4 (a) @(46,29) /sn:0 /w:[ 0 ]
  //: OUT g3 (cout) @(268,143) /sn:0 /w:[ 0 ]
  exor g2 (.b(b), .a(a), .cout(s));   //: @(96, 18) /sz:(99, 55) /sn:0 /p:[ Li0>0 Li1>3 Ro0<1 ]
  //: OUT g1 (s) @(268,41) /sn:0 /w:[ 0 ]
  //: joint g6 (b) @(65, 156) /w:[ 2 1 4 -1 ]
  //: joint g7 (a) @(79, 29) /w:[ 2 1 -1 4 ]
  //: IN g5 (b) @(50,156) /sn:0 /w:[ 5 ]
  and0 g0 (.a(a), .b(b), .cout(cout));   //: @(166, 120) /sz:(77, 48) /sn:0 /p:[ Li0>5 Li1>3 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin full_adder
module full_adder(b, a, s, cout, cin);
//: interface  /sz:(57, 74) /bd:[ Ti0>a(13/57) Ti1>b(42/57) Ri0>cin(50/74) Lo0<cout(48/74) Bo0<s(28/57) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(127,51)(127,107)(127,107)(127,84){1}
input cin;    //: /sn:0 {0}(39,172)(134,172)(134,219){1}
output s;    //: /sn:0 {0}(97,294)(97,295)(97,295)(97,330){1}
input a;    //: /sn:0 {0}(83,50)(83,106)(83,106)(83,84){1}
output cout;    //: /sn:0 {0}(272,274)(262,274)(262,274)(297,274){1}
wire w0;    //: /sn:0 {0}(90,159)(90,216)(90,216)(90,219){1}
wire w1;    //: /sn:0 {0}(191,277)(188,277)(188,277)(213,277){1}
wire w2;    //: /sn:0 {0}(184,142)(201,142)(201,249)(213,249){1}
//: enddecls

  //: IN g4 (b) @(127,49) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (a) @(83,48) /sn:0 /R:3 /w:[ 0 ]
  or0 g2 (.a(w2), .b(w1), .cout(cout));   //: @(214, 240) /sz:(57, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  half_adder g1 (.a(w0), .b(cin), .s(s), .cout(w1));   //: @(67, 220) /sz:(123, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Ro0<0 ]
  //: OUT g6 (s) @(97,327) /sn:0 /R:3 /w:[ 1 ]
  //: OUT g7 (cout) @(294,274) /sn:0 /w:[ 1 ]
  //: IN g5 (cin) @(37,172) /sn:0 /w:[ 0 ]
  half_adder g0 (.a(a), .b(b), .s(w0), .cout(w2));   //: @(60, 85) /sz:(123, 73) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Ro0<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin complemento
module complemento(cout, b);
//: interface  /sz:(194, 51) /bd:[ Ti0>b[3:0](95/194) Bo0<cout[3:0](100/194) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:491,146)(413,146){1}
//: {2}(412,146)(334,146){3}
//: {4}(333,146)(261,146){5}
//: {6}(260,146)(185,146){7}
//: {8}(184,146)(#:147,146){9}
supply1 w4;    //: /sn:0 {0}(328,65)(328,86){1}
//: {2}(330,88)(360,88){3}
//: {4}(364,88)(441,88)(441,178){5}
//: {6}(362,90)(362,178){7}
//: {8}(326,88)(291,88){9}
//: {10}(287,88)(213,88)(213,178){11}
//: {12}(289,90)(289,179){13}
output [3:0] cout;    //: /sn:0 {0}(313,457)(#:313,388){1}
wire w6;    //: /sn:0 {0}(334,150)(334,178){1}
wire w3;    //: /sn:0 {0}(261,179)(261,150){1}
wire w0;    //: /sn:0 {0}(185,150)(185,178){1}
wire w8;    //: /sn:0 {0}(318,382)(318,353)(350,353)(350,279){1}
wire w11;    //: /sn:0 {0}(429,279)(429,365)(328,365)(328,382){1}
wire w2;    //: /sn:0 {0}(201,279)(201,367)(298,367)(298,382){1}
wire w5;    //: /sn:0 {0}(308,382)(308,353)(277,353)(277,280){1}
wire w9;    //: /sn:0 {0}(413,150)(413,178){1}
//: enddecls

  assign w6 = b[2]; //: TAP g8 @(334,144) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  exor g4 (.a(w4), .b(w9), .cout(w11));   //: @(398, 179) /sz:(55, 99) /R:3 /sn:0 /p:[ Ti0>5 Ti1>1 Bo0<0 ]
  //: joint g13 (w4) @(362, 88) /w:[ 4 -1 3 6 ]
  exor g3 (.a(w4), .b(w6), .cout(w8));   //: @(319, 179) /sz:(55, 99) /R:3 /sn:0 /p:[ Ti0>7 Ti1>1 Bo0<1 ]
  exor g2 (.a(w4), .b(w3), .cout(w5));   //: @(246, 180) /sz:(55, 99) /R:3 /sn:0 /p:[ Ti0>13 Ti1>0 Bo0<1 ]
  exor g1 (.a(w4), .b(w0), .cout(w2));   //: @(170, 179) /sz:(55, 99) /R:3 /sn:0 /p:[ Ti0>11 Ti1>1 Bo0<0 ]
  assign w9 = b[3]; //: TAP g11 @(413,144) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  assign w0 = b[0]; //: TAP g6 @(185,144) /sn:0 /R:1 /w:[ 0 8 7 ] /ss:1
  assign w3 = b[1]; //: TAP g7 @(261,144) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  //: OUT g9 (cout) @(313,454) /sn:0 /R:3 /w:[ 0 ]
  //: joint g15 (w4) @(328, 88) /w:[ 2 1 8 -1 ]
  assign cout = {w11, w8, w5, w2}; //: CONCAT g5  @(313,387) /sn:0 /R:3 /w:[ 1 1 0 0 1 ] /dr:0 /tp:0 /drp:1
  //: VDD g14 (w4) @(339,65) /sn:0 /w:[ 0 ]
  //: IN g0 (b) @(145,146) /sn:0 /w:[ 9 ]
  //: joint g12 (w4) @(289, 88) /w:[ 9 -1 10 12 ]

endmodule
//: /netlistEnd

//: /netlistBegin inverter
module inverter(a, cout);
//: interface  /sz:(123, 48) /bd:[ Li0>a(23/48) Ro0<cout(21/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w0;    //: /sn:0 {0}(235,243)(235,233)(235,233)(235,199){1}
supply0 w1;    //: /sn:0 {0}(235,383)(235,337){1}
input a;    //: /sn:0 {0}(122,288)(188,288){1}
//: {2}(190,286)(190,251)(221,251){3}
//: {4}(190,290)(190,328)(221,328){5}
output cout;    //: /sn:0 {0}(235,320)(235,289){1}
//: {2}(237,287)(306,287)(306,288)(308,288){3}
//: {4}(235,285)(235,271)(235,271)(235,260){5}
//: enddecls

  //: IN g4 (a) @(120,288) /sn:0 /w:[ 0 ]
  _GGNMOS #(2, 1) g3 (.Z(cout), .S(w1), .G(a));   //: @(229,328) /sn:0 /w:[ 0 1 5 ]
  _GGPMOS #(2, 1) g2 (.Z(cout), .S(w0), .G(a));   //: @(229,251) /sn:0 /w:[ 5 0 3 ]
  //: GROUND g1 (w1) @(235,389) /sn:0 /w:[ 0 ]
  //: OUT g6 (cout) @(305,288) /sn:0 /w:[ 3 ]
  //: joint g7 (cout) @(235, 287) /w:[ 2 4 -1 1 ]
  //: joint g5 (a) @(190, 288) /w:[ -1 2 1 4 ]
  //: VDD g0 (w0) @(246,199) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin shift1
module shift1(s, cout, bit_succ, a);
//: interface  /sz:(100, 122) /bd:[ Ti0>a(76/100) Ti1>bit_succ(30/100) Li0>s(27/122) Bo0<cout(51/100) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input bit_succ;    //: /sn:0 {0}(309,154)(309,68)(262,68)(262,-65){1}
input s;    //: /sn:0 {0}(153,-21)(335,-21){1}
//: {2}(339,-21)(420,-21)(420,-11){3}
//: {4}(337,-19)(337,154){5}
input a;    //: /sn:0 {0}(370,-62)(370,142)(394,142)(394,154){1}
output cout;    //: /sn:0 {0}(352,347)(352,407){1}
wire w4;    //: /sn:0 {0}(422,114)(422,154){1}
wire w2;    //: /sn:0 {0}(322,233)(322,273)(349,273)(349,288){1}
wire w5;    //: /sn:0 {0}(407,233)(407,275)(377,275)(377,288){1}
//: enddecls

  //: IN g8 (s) @(151,-21) /sn:0 /w:[ 0 ]
  //: OUT g4 (cout) @(352,404) /sn:0 /R:3 /w:[ 1 ]
  or0 g3 (.a(w5), .b(w2), .cout(cout));   //: @(338, 289) /sz:(48, 57) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]
  and0 g2 (.a(w4), .b(a), .cout(w5));   //: @(382, 155) /sz:(48, 77) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 ]
  and0 g1 (.a(s), .b(bit_succ), .cout(w2));   //: @(297, 155) /sz:(48, 77) /R:3 /sn:0 /p:[ Ti0>5 Ti1>0 Bo0<0 ]
  //: joint g6 (s) @(337, -21) /w:[ 2 -1 1 4 ]
  //: IN g7 (bit_succ) @(262,-67) /sn:0 /R:3 /w:[ 1 ]
  inverter g5 (.a(s), .cout(w4));   //: @(395, -10) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>3 Bo0<0 ]
  //: IN g0 (a) @(370,-64) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin or4
module or4(d, c, b, cout, a);
//: interface  /sz:(73, 79) /bd:[ Ti0>a(15/73) Ti1>b(32/73) Ti2>c(45/73) Ti3>d(63/73) Bo0<cout(39/73) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(308,173)(328,173)(328,173)(350,173){1}
input d;    //: /sn:0 {0}(351,227)(330,227)(330,227)(308,227){1}
input a;    //: /sn:0 {0}(308,145)(327,145)(327,145)(350,145){1}
output cout;    //: /sn:0 {0}(523,212)(558,212){1}
input c;    //: /sn:0 {0}(351,199)(329,199)(329,199)(308,199){1}
wire w2;    //: /sn:0 {0}(409,170)(426,170)(426,187)(464,187){1}
wire w5;    //: /sn:0 {0}(464,215)(425,215)(425,224)(410,224){1}
//: enddecls

  or0 g4 (.b(b), .a(a), .cout(w2));   //: @(351, 136) /sz:(57, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g3 (d) @(306,227) /sn:0 /w:[ 1 ]
  //: IN g2 (c) @(306,199) /sn:0 /w:[ 1 ]
  //: IN g1 (b) @(306,173) /sn:0 /w:[ 0 ]
  or0 g6 (.b(w5), .a(w2), .cout(cout));   //: @(465, 178) /sz:(57, 48) /sn:0 /p:[ Li0>0 Li1>1 Ro0<0 ]
  //: OUT g7 (cout) @(555,212) /sn:0 /w:[ 1 ]
  or0 g5 (.b(d), .a(c), .cout(w5));   //: @(352, 190) /sz:(57, 48) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: IN g0 (a) @(306,145) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin and4
module and4(d, c, b, cout, a);
//: interface  /sz:(82, 82) /bd:[ Li0>d(71/82) Li1>c(54/82) Li2>b(36/82) Li3>a(17/82) Ro0<cout(48/82) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(321,178)(272,178){1}
input d;    //: /sn:0 {0}(321,235)(275,235){1}
input a;    //: /sn:0 {0}(321,150)(270,150){1}
output cout;    //: /sn:0 {0}(573,193)(537,193){1}
input c;    //: /sn:0 {0}(321,207)(272,207){1}
wire w2;    //: /sn:0 {0}(458,178)(415,178)(415,165)(400,165){1}
wire w5;    //: /sn:0 {0}(458,206)(415,206)(415,222)(400,222){1}
//: enddecls

  and0 g4 (.a(a), .b(b), .cout(w2));   //: @(322, 142) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: IN g3 (d) @(273,235) /sn:0 /w:[ 1 ]
  //: IN g2 (c) @(270,207) /sn:0 /w:[ 1 ]
  //: IN g1 (b) @(270,178) /sn:0 /w:[ 1 ]
  and0 g6 (.a(w2), .b(w5), .cout(cout));   //: @(459, 170) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: OUT g7 (cout) @(570,193) /sn:0 /w:[ 0 ]
  and0 g5 (.a(c), .b(d), .cout(w5));   //: @(322, 199) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  //: IN g0 (a) @(268,150) /sn:0 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin mux4
module mux4(a, s, b, cout);
//: interface  /sz:(127, 40) /bd:[ Ti0>a[3:0](37/127) Ti1>b[3:0](88/127) Li0>s(24/40) Ro0<cout[3:0](23/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:68,31)(68,91){1}
//: {2}(68,92)(68,175){3}
//: {4}(68,176)(68,282){5}
//: {6}(68,283)(68,365){7}
//: {8}(68,366)(68,388){9}
input s;    //: /sn:0 {0}(102,78)(102,133){1}
//: {2}(104,135)(132,135){3}
//: {4}(102,137)(102,227){5}
//: {6}(104,229)(128,229){7}
//: {8}(102,231)(102,331){9}
//: {10}(104,333)(128,333){11}
//: {12}(102,335)(102,432)(129,432){13}
input [3:0] a;    //: /sn:0 {0}(#:42,32)(42,97){1}
//: {2}(42,98)(42,187){3}
//: {4}(42,188)(42,293){5}
//: {6}(42,294)(42,370){7}
//: {8}(42,371)(42,391){9}
output [3:0] cout;    //: /sn:0 {0}(#:369,261)(412,261){1}
wire w7;    //: /sn:0 {0}(363,266)(329,266)(329,330)(235,330){1}
wire w15;    //: /sn:0 {0}(236,429)(349,429)(349,276)(363,276){1}
wire w4;    //: /sn:0 {0}(72,283)(197,283)(197,312){1}
wire w3;    //: /sn:0 {0}(363,256)(329,256)(329,226)(235,226){1}
wire w0;    //: /sn:0 {0}(72,176)(197,176)(197,208){1}
wire w1;    //: /sn:0 {0}(46,188)(160,188)(160,208){1}
wire w8;    //: /sn:0 {0}(72,92)(201,92)(201,114){1}
wire w12;    //: /sn:0 {0}(72,366)(198,366)(198,411){1}
wire w11;    //: /sn:0 {0}(239,132)(348,132)(348,246)(363,246){1}
wire w13;    //: /sn:0 {0}(46,371)(161,371)(161,411){1}
wire w5;    //: /sn:0 {0}(46,294)(160,294)(160,312){1}
wire w9;    //: /sn:0 {0}(46,98)(164,98)(164,114){1}
//: enddecls

  //: IN g8 (a) @(42,30) /sn:0 /R:3 /w:[ 0 ]
  //: IN g4 (s) @(102,76) /sn:0 /R:3 /w:[ 0 ]
  assign w13 = a[3]; //: TAP g13 @(40,371) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  mux1 g3 (.a(w13), .b(w12), .s(s), .cout(w15));   //: @(130, 412) /sz:(105, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>13 Ro0<0 ]
  mux1 g2 (.a(w9), .b(w8), .s(s), .cout(w11));   //: @(133, 115) /sz:(105, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>3 Ro0<0 ]
  mux1 g1 (.a(w5), .b(w4), .s(s), .cout(w7));   //: @(129, 313) /sz:(105, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>11 Ro0<1 ]
  assign w0 = b[1]; //: TAP g16 @(66,176) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  assign w1 = a[1]; //: TAP g11 @(40,188) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  assign w9 = a[0]; //: TAP g10 @(40,98) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  assign cout = {w15, w7, w3, w11}; //: CONCAT g19  @(368,261) /sn:0 /w:[ 0 1 0 0 1 ] /dr:1 /tp:0 /drp:1
  //: joint g6 (s) @(102, 229) /w:[ 6 5 -1 8 ]
  //: IN g9 (b) @(68,29) /sn:0 /R:3 /w:[ 0 ]
  //: joint g7 (s) @(102, 333) /w:[ 10 9 -1 12 ]
  assign w4 = b[2]; //: TAP g15 @(66,283) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  assign w8 = b[0]; //: TAP g17 @(66,92) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  assign w12 = b[3]; //: TAP g14 @(66,366) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: joint g5 (s) @(102, 135) /w:[ 2 1 -1 4 ]
  mux1 g0 (.a(w1), .b(w0), .s(s), .cout(w3));   //: @(129, 209) /sz:(105, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>7 Ro0<1 ]
  //: OUT g18 (cout) @(409,261) /sn:0 /w:[ 1 ]
  assign w5 = a[2]; //: TAP g12 @(40,294) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin nor0
module nor0(cout, a, b);
//: interface  /sz:(62, 50) /bd:[ Li0>a(9/50) Li1>b(39/50) Ro0<cout(34/50) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(137,370)(224,370)(224,370)(189,370){1}
//: {2}(193,370)(274,370)(274,370)(323,370){3}
//: {4}(191,368)(191,222)(251,222){5}
supply1 w4;    //: /sn:0 {0}(265,105)(265,155){1}
supply0 w1;    //: /sn:0 {0}(279,448)(279,414){1}
//: {2}(281,412)(337,412)(337,379){3}
//: {4}(277,412)(214,412)(214,328){5}
input a;    //: /sn:0 {0}(137,163)(200,163)(200,163)(157,163){1}
//: {2}(161,163)(222,163)(222,163)(251,163){3}
//: {4}(159,165)(159,319)(200,319){5}
output cout;    //: /sn:0 {0}(214,311)(214,283)(263,283){1}
//: {2}(267,283)(337,283)(337,362){3}
//: {4}(265,281)(265,250){5}
//: {6}(267,248)(296,248)(296,248)(342,248){7}
//: {8}(265,246)(265,231){9}
wire w0;    //: /sn:0 {0}(265,214)(265,172){1}
//: enddecls

  //: OUT g4 (cout) @(339,248) /sn:0 /w:[ 7 ]
  //: joint g8 (cout) @(265, 283) /w:[ 2 4 1 -1 ]
  //: IN g3 (a) @(135,163) /sn:0 /w:[ 0 ]
  //: joint g13 (b) @(191, 370) /w:[ 2 4 1 -1 ]
  //: VDD g2 (w4) @(276,105) /sn:0 /w:[ 0 ]
  _GGPMOS #(2, 1) g1 (.Z(cout), .S(w0), .G(b));   //: @(259,222) /sn:0 /w:[ 9 0 5 ]
  //: IN g11 (b) @(135,370) /sn:0 /w:[ 0 ]
  //: joint g10 (w1) @(279, 412) /w:[ 2 -1 4 1 ]
  _GGNMOS #(2, 1) g6 (.Z(cout), .S(w1), .G(a));   //: @(208,319) /sn:0 /w:[ 0 5 5 ]
  _GGNMOS #(2, 1) g7 (.Z(cout), .S(w1), .G(b));   //: @(331,370) /sn:0 /w:[ 3 3 3 ]
  //: GROUND g9 (w1) @(279,454) /sn:0 /w:[ 0 ]
  //: joint g5 (cout) @(265, 248) /w:[ 6 8 -1 5 ]
  _GGPMOS #(2, 1) g0 (.Z(w0), .S(w4), .G(a));   //: @(259,163) /sn:0 /w:[ 1 1 3 ]
  //: joint g12 (a) @(159, 163) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin comparatore1
module comparatore1(b, magg, equal, a, minor);
//: interface  /sz:(110, 122) /bd:[ Ti0>b(74/110) Ti1>a(20/110) Bo0<minor(76/110) Bo1<magg(25/110) Ro0<equal(101/122) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(340,387)(236,387)(236,320){1}
//: {2}(238,318)(249,318)(249,224)(335,224){3}
//: {4}(234,318)(69,318){5}
//: {6}(65,318)(40,318){7}
//: {8}(67,320)(67,357)(93,357){9}
output equal;    //: /sn:0 {0}(549,265)(634,265){1}
output minor;    //: /sn:0 {0}(419,374)(635,374){1}
output magg;    //: /sn:0 {0}(413,134)(635,134){1}
input a;    //: /sn:0 {0}(335,196)(248,196)(248,121){1}
//: {2}(250,119)(334,119){3}
//: {4}(246,119)(79,119){5}
//: {6}(75,119)(58,119){7}
//: {8}(77,121)(77,176)(93,176){9}
wire w4;    //: /sn:0 {0}(340,359)(266,359)(266,176){1}
//: {2}(268,174)(321,174)(321,281)(335,281){3}
//: {4}(264,174)(218,174){5}
wire w3;    //: /sn:0 {0}(335,309)(289,309){1}
//: {2}(287,307)(287,147)(334,147){3}
//: {4}(287,311)(287,355)(218,355){5}
wire w2;    //: /sn:0 {0}(414,211)(475,211)(475,240)(490,240){1}
wire w5;    //: /sn:0 {0}(414,296)(475,296)(475,268)(490,268){1}
//: enddecls

  or0 g4 (.a(w2), .b(w5), .cout(equal));   //: @(491, 231) /sz:(57, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: IN g8 (b) @(38,318) /sn:0 /w:[ 7 ]
  and0 g3 (.a(w4), .b(b), .cout(minor));   //: @(341, 351) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>0 Ro0<0 ]
  //: joint g13 (a) @(77, 119) /w:[ 5 -1 6 8 ]
  and0 g2 (.a(a), .b(w3), .cout(magg));   //: @(335, 111) /sz:(77, 48) /sn:0 /p:[ Li0>3 Li1>3 Ro0<0 ]
  and0 g1 (.a(w4), .b(w3), .cout(w5));   //: @(336, 273) /sz:(77, 48) /sn:0 /p:[ Li0>3 Li1>0 Ro0<0 ]
  //: OUT g11 (magg) @(632,134) /sn:0 /w:[ 1 ]
  //: joint g16 (b) @(236, 318) /w:[ 2 -1 4 1 ]
  //: OUT g10 (equal) @(631,265) /sn:0 /w:[ 1 ]
  inverter g6 (.a(a), .cout(w4));   //: @(94, 153) /sz:(123, 48) /sn:0 /p:[ Li0>9 Ro0<5 ]
  //: IN g7 (a) @(56,119) /sn:0 /w:[ 7 ]
  //: OUT g9 (minor) @(632,374) /sn:0 /w:[ 1 ]
  //: joint g15 (w3) @(287, 309) /w:[ 1 2 -1 4 ]
  //: joint g17 (w4) @(266, 174) /w:[ 2 -1 4 1 ]
  inverter g5 (.a(b), .cout(w3));   //: @(94, 334) /sz:(123, 48) /sn:0 /p:[ Li0>9 Ro0<5 ]
  //: joint g14 (a) @(248, 119) /w:[ 2 -1 4 1 ]
  and0 g0 (.a(a), .b(b), .cout(w2));   //: @(336, 188) /sz:(77, 48) /sn:0 /p:[ Li0>0 Li1>3 Ro0<0 ]
  //: joint g12 (b) @(67, 318) /w:[ 5 -1 6 8 ]

endmodule
//: /netlistEnd

//: /netlistBegin mux1
module mux1(cout, a, b, s);
//: interface  /sz:(105, 40) /bd:[ Ti0>b(68/105) Ti1>a(31/105) Li0>s(20/40) Ro0<cout(17/40) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input b;    //: /sn:0 {0}(310,352)(264,352){1}
input s;    //: /sn:0 {0}(190,108)(190,124){1}
//: {2}(192,126)(221,126)(221,137){3}
//: {4}(190,128)(190,380)(310,380){5}
input a;    //: /sn:0 {0}(310,289)(275,289)(275,290)(260,290){1}
output cout;    //: /sn:0 {0}(493,349)(550,349){1}
wire w6;    //: /sn:0 {0}(389,367)(419,367)(419,352)(434,352){1}
wire w0;    //: /sn:0 {0}(223,262)(223,315)(235,315)(235,317)(310,317){1}
wire w3;    //: /sn:0 {0}(389,304)(419,304)(419,324)(434,324){1}
//: enddecls

  //: OUT g8 (cout) @(547,349) /sn:0 /w:[ 1 ]
  and0 g4 (.b(s), .a(b), .cout(w6));   //: @(311, 344) /sz:(77, 48) /sn:0 /p:[ Li0>5 Li1>0 Ro0<0 ]
  and0 g3 (.b(w0), .a(a), .cout(w3));   //: @(311, 281) /sz:(77, 48) /sn:0 /p:[ Li0>1 Li1>0 Ro0<0 ]
  //: IN g2 (a) @(258,290) /sn:0 /w:[ 1 ]
  inverter g1 (.a(s), .cout(w0));   //: @(196, 138) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>3 Bo0<0 ]
  or0 g6 (.b(w6), .a(w3), .cout(cout));   //: @(435, 315) /sz:(57, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<0 ]
  //: joint g7 (s) @(190, 126) /w:[ 2 1 -1 4 ]
  //: IN g5 (b) @(262,352) /sn:0 /w:[ 1 ]
  //: IN g0 (s) @(190,106) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin exor
module exor(b, a, cout);
//: interface  /sz:(99, 55) /bd:[ Li0>b(39/55) Li1>a(11/55) Ro0<cout(23/55) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(136,287)(152,287)(152,287)(160,287){1}
//: {2}(164,287)(342,287){3}
//: {4}(162,285)(162,169)(192,169){5}
input a;    //: /sn:0 {0}(194,246)(176,246)(176,138){1}
//: {2}(176,134)(176,124)(316,124)(316,124)(345,124){3}
//: {4}(174,136)(167,136)(167,136)(136,136){5}
output cout;    //: /sn:0 {0}(587,211)(561,211){1}
wire w6;    //: /sn:0 {0}(466,187)(453,187)(453,148)(440,148){1}
wire w7;    //: /sn:0 {0}(466,230)(456,230)(456,268)(437,268){1}
wire w4;    //: /sn:0 {0}(345,167)(317,167){1}
wire w3;    //: /sn:0 {0}(342,244)(319,244){1}
//: enddecls

  //: IN g4 (b) @(134,287) /sn:0 /w:[ 0 ]
  nand0 g8 (.b(w7), .a(w6), .cout(cout));   //: @(467, 176) /sz:(93, 70) /sn:0 /p:[ Li0>0 Li1>0 Ro0<1 ]
  inverter g3 (.a(a), .cout(w3));   //: @(195, 223) /sz:(123, 48) /sn:0 /p:[ Li0>0 Ro0<1 ]
  inverter g2 (.a(b), .cout(w4));   //: @(193, 146) /sz:(123, 48) /sn:0 /p:[ Li0>5 Ro0<1 ]
  //: IN g1 (a) @(134,136) /sn:0 /w:[ 5 ]
  //: joint g6 (a) @(176, 136) /w:[ -1 2 4 1 ]
  //: OUT g9 (cout) @(584,211) /sn:0 /w:[ 0 ]
  //: joint g7 (b) @(162, 287) /w:[ 2 4 1 -1 ]
  nand0 g5 (.b(b), .a(w3), .cout(w7));   //: @(343, 233) /sz:(93, 70) /sn:0 /p:[ Li0>3 Li1>0 Ro0<1 ]
  nand0 g0 (.b(w4), .a(a), .cout(w6));   //: @(346, 113) /sz:(93, 70) /sn:0 /p:[ Li0>0 Li1>3 Ro0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin comparatore4
module comparatore4(b, a, c);
//: interface  /sz:(181, 114) /bd:[ Li0>a[3:0](24/114) Li1>b[3:0](77/114) Ro0<c(54/114) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input [3:0] b;    //: /sn:0 {0}(#:82,215)(201,215){1}
//: {2}(202,215)(347,215){3}
//: {4}(348,215)(500,215){5}
//: {6}(501,215)(671,215){7}
//: {8}(672,215)(682,215){9}
input [3:0] a;    //: /sn:0 {0}(#:82,166)(147,166){1}
//: {2}(148,166)(293,166){3}
//: {4}(294,166)(446,166){5}
//: {6}(447,166)(617,166){7}
//: {8}(618,166)(635,166){9}
output c;    //: /sn:0 {0}(351,868)(351,814){1}
wire w6;    //: /sn:0 {0}(348,219)(348,265){1}
wire w7;    //: /sn:0 {0}(600,600)(600,570)(623,570)(623,391){1}
wire w16;    //: /sn:0 {0}(503,390)(503,412)(509,412)(509,417){1}
wire w14;    //: /sn:0 {0}(452,390)(452,554)(436,554)(436,593){1}
wire w4;    //: /sn:0 {0}(166,661)(166,718)(327,718)(327,733){1}
wire w15;    //: /sn:0 {0}(248,583)(248,568){1}
//: {2}(250,566)(401,566)(401,581){3}
//: {4}(403,583)(546,583)(546,600){5}
//: {6}(401,585)(401,593){7}
//: {8}(248,564)(248,529)(256,529)(256,369)(239,369){9}
wire w3;    //: /sn:0 {0}(153,391)(153,489)(153,489)(153,582){1}
wire w0;    //: /sn:0 {0}(148,170)(148,267){1}
wire w34;    //: /sn:0 {0}(278,583)(278,552)(359,552)(359,542){1}
wire w21;    //: /sn:0 {0}(663,417)(663,401)(674,401)(674,391){1}
wire w43;    //: /sn:0 {0}(665,542)(665,573)(653,573)(653,591)(619,591)(619,600){1}
wire w28;    //: /sn:0 {0}(385,367)(418,367)(418,566){1}
//: {2}(420,568)(563,568)(563,600){3}
//: {4}(418,570)(418,593){5}
wire w23;    //: /sn:0 {0}(511,542)(511,578)(455,578)(455,593){1}
wire w41;    //: /sn:0 {0}(181,582)(181,557)(200,557)(200,542){1}
wire w24;    //: /sn:0 {0}(344,733)(344,699)(262,699)(262,660){1}
wire w36;    //: /sn:0 {0}(583,698)(583,718)(375,718)(375,733){1}
wire w1;    //: /sn:0 {0}(202,219)(202,267){1}
wire w8;    //: /sn:0 {0}(263,583)(263,538)(299,538)(299,389){1}
wire w18;    //: /sn:0 {0}(583,600)(583,368)(538,368){1}
wire w12;    //: /sn:0 {0}(618,170)(618,267){1}
wire w11;    //: /sn:0 {0}(501,219)(501,266){1}
wire w2;    //: /sn:0 {0}(718,369)(709,369){1}
wire w10;    //: /sn:0 {0}(447,170)(447,266){1}
wire w13;    //: /sn:0 {0}(672,219)(672,267){1}
wire w27;    //: /sn:0 {0}(357,733)(357,692)(424,692)(424,677){1}
wire w5;    //: /sn:0 {0}(294,170)(294,265){1}
wire w9;    //: /sn:0 {0}(350,389)(350,411)(357,411)(357,417){1}
wire w42;    //: /sn:0 {0}(204,391)(204,407)(198,407)(198,417){1}
//: enddecls

  assign w5 = a[2]; //: TAP g8 @(294,164) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w0 = a[3]; //: TAP g4 @(148,164) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w11 = b[1]; //: TAP g13 @(501,213) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w1 = b[3]; //: TAP g3 @(202,213) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  comparatore1 g2 (.b(w1), .a(w0), .minor(w42), .magg(w3), .equal(w15));   //: @(128, 268) /sz:(110, 122) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 Ro0<9 ]
  //: IN g1 (b) @(80,215) /sn:0 /w:[ 0 ]
  inverter g16 (.a(w16), .cout(w23));   //: @(484, 418) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>1 Bo0<0 ]
  comparatore1 g11 (.b(w13), .a(w12), .minor(w21), .magg(w7), .equal(w2));   //: @(598, 268) /sz:(110, 122) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Bo1<1 Ro0<1 ]
  comparatore1 g10 (.b(w11), .a(w10), .minor(w16), .magg(w14), .equal(w18));   //: @(427, 267) /sz:(110, 122) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 Ro0<1 ]
  and3 g19 (.c(w15), .b(w8), .a(w34), .cout(w24));   //: @(235, 584) /sz:(57, 75) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Bo0<1 ]
  inverter g6 (.a(w42), .cout(w41));   //: @(173, 418) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>1 Bo0<1 ]
  inverter g7 (.a(w9), .cout(w34));   //: @(332, 418) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>1 Bo0<1 ]
  assign w6 = b[2]; //: TAP g9 @(348,213) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w13 = b[0]; //: TAP g15 @(672,213) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  and4 g20 (.d(w15), .c(w28), .b(w14), .a(w23), .cout(w27));   //: @(390, 594) /sz:(82, 82) /R:3 /sn:0 /p:[ Ti0>7 Ti1>5 Ti2>1 Ti3>1 Bo0<1 ]
  or4 g25 (.d(w36), .c(w27), .b(w24), .a(w4), .cout(c));   //: @(312, 734) /sz:(73, 79) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Ti3>1 Bo0<1 ]
  inverter g17 (.a(w21), .cout(w43));   //: @(638, 418) /sz:(48, 123) /R:3 /sn:0 /p:[ Ti0>0 Bo0<0 ]
  assign w12 = a[0]; //: TAP g14 @(618,164) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  comparatore1 g5 (.b(w6), .a(w5), .minor(w9), .magg(w8), .equal(w28));   //: @(274, 266) /sz:(110, 122) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<1 Ro0<0 ]
  and5 g21 (.e(w15), .d(w28), .c(w18), .b(w7), .a(w43), .cout(w36));   //: @(533, 601) /sz:(94, 96) /R:3 /sn:0 /p:[ Ti0>5 Ti1>3 Ti2>0 Ti3>0 Ti4>1 Bo0<0 ]
  //: joint g24 (w15) @(401, 583) /w:[ 4 3 -1 6 ]
  //: joint g23 (w28) @(418, 568) /w:[ 2 1 -1 4 ]
  //: IN g0 (a) @(80,166) /sn:0 /w:[ 0 ]
  //: joint g22 (w15) @(248, 566) /w:[ 2 8 -1 1 ]
  and0 g18 (.b(w3), .a(w41), .cout(w4));   //: @(141, 583) /sz:(48, 77) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Bo0<0 ]
  assign w10 = a[1]; //: TAP g12 @(447,164) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: OUT g33 (c) @(351,865) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

